//register ex/mem
`timescale 1ns/1ps
`include "defines.v"

module r_ex_mem(
    
);

endmodule